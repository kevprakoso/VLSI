module scaler(
input wire [23:0] data_in,
input wire [4:0] step
output reg [23:0] data_out
)