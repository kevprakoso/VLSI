module  calc (  
	angle_in,
	count_n,
	mag,
	right_p,
	left_p
	);
	
input		angle_in;
input		count_n;
input		mag;
output	right_p;
output	left_p;

endmodule