module  adjust (  
	angle_in,
	angle_out,
	count_n
	);
	
input		angle_in;
output		angle_out;
output		count_n;

endmodule
