


module calculateScaleStep(
	rows,
	cols
	step
);

input	rows;
input	cols;
output  [5:0] step;




