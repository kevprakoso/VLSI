module histogram (  
	count_n,
	right_p,
	left_p,
	output_h
	);
	
input		count_n;
input	right_p;
input	left_p;
output output_h;

endmodule